module servo_pos_dcd (
    input  wire [ 7:0] deg,

    output wire [19:0] pos
);

    /* decode degrees (0-180) to servo PMW bound */

endmodule
